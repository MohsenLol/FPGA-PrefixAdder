module BrentKung64b (A, B, S);
input [63 : 0] A;
input [63 : 0] B;
output [64 : 0] S;
wire g_2_0_61, c [64 : 0], g_2_0_29, p_4_16_31, g_1_34_35, g_0_25_25, p_0_26_26, g_1_0_44, p_0_47_47, p_0_18_18, g_2_60_63, p_1_34_35, p_1_46_47, p_0_46_46, p_0_4_4, g_0_21_21, g_3_0_51, g_1_0_22, p_0_61_61, p_2_16_19, p_0_60_60, g_0_51_51, p_3_56_63, g_1_44_45, p_1_12_13, g_1_0_62, g_1_32_33, g_1_0_56, p_1_16_17, p_0_9_9, g_2_0_45, g_0_17_17, g_1_54_55, g_1_0_38, p_0_21_21, g_0_30_30, g_0_15_15, g_1_42_43, g_4_32_47, g_0_57_57, g_0_43_43, g_1_0_20, g_4_0_23, p_0_8_8, p_0_48_48, p_3_16_23, g_0_9_9, p_1_40_41, g_1_38_39, g_1_22_23, g_0_42_42, p_0_17_17, p_0_2_2, p_0_10_10, g_0_7_7, g_0_32_32, g_1_4_5, g_3_0_59, g_0_3_3, g_1_26_27, g_1_0_6, g_0_26_26, g_2_52_55, g_0_1_1, g_3_56_63, p_1_22_23, g_1_60_61, p_4_48_63, p_1_60_61, g_0_37_37, p_0_30_30, p_1_62_63, g_1_30_31, g_0_14_14, g_1_0_10, p_0_5_5, g_3_40_47, g_2_0_53, g_0_56_56, g_2_0_41, p_2_48_51, p_1_2_3, p_1_14_15, g_0_19_19, g_1_58_59, g_2_16_19, g_0_38_38, g_1_40_41, p_1_58_59, g_0_61_61, g_1_0_58, g_2_32_35, g_4_48_63, g_0_8_8, g_1_12_13, g_1_0_36, g_1_50_51, p_0_41_41, g_1_0_8, p_0_15_15, p_0_31_31, g_3_24_31, g_4_0_15, p_2_60_63, p_2_28_31, p_0_13_13, p_0_25_25, p_0_51_51, g_3_0_19, p_2_36_39, g_1_0_52, g_1_0_26, g_1_6_7, p_1_50_51, g_1_36_37, g_3_16_23, g_2_48_51, g_1_0_50, g_2_44_47, p_0_3_3, p_1_6_7, p_1_44_45, p_0_6_6, g_0_63_63, p_0_0_0, p_0_52_52, g_0_40_40, g_0_10_10, g_2_0_17, p_0_58_58, g_0_28_28, g_2_0_5, p_1_56_57, g_0_54_54, g_0_52_52, g_0_24_24, g_0_16_16, p_1_38_39, g_1_56_57, p_1_32_33, g_1_0_34, p_0_28_28, g_0_58_58, p_0_55_55, p_0_42_42, g_0_47_47, g_3_48_55, g_1_0_46, p_1_8_9, p_0_14_14, g_2_28_31, g_0_20_20, p_1_52_53, p_4_32_47, g_0_35_35, g_3_0_11, g_1_0_54, p_2_12_15, g_1_0_42, g_3_0_35, p_3_24_31, g_5_32_63, g_0_2_2, g_1_28_29, p_2_40_43, p_0_62_62, g_2_0_13, g_0_22_22, g_0_11_11, g_0_23_23, g_0_46_46, p_2_24_27, g_2_0_3, g_0_60_60, p_5_32_63, p_0_29_29, g_1_0_12, p_1_28_29, g_0_59_59, g_0_41_41, g_0_34_34, p_1_24_25, g_1_0_1, p_0_36_36, p_2_56_59, g_0_50_50, p_1_18_19, g_2_56_59, p_3_8_15, g_1_10_11, p_0_19_19, p_0_44_44, g_1_48_49, g_2_8_11, p_0_40_40, p_3_48_55, g_0_29_29, g_2_0_49, g_1_18_19, g_3_0_7, p_0_7_7, g_0_6_6, g_0_0_0, p_3_32_39, p_0_22_22, g_1_8_9, g_2_40_43, p_0_38_38, p_0_63_63, p_2_8_11, g_1_0_16, p_0_37_37, p_0_27_27, p_0_35_35, p_2_52_55, g_2_36_39, p_0_49_49, g_1_0_32, g_2_12_15, g_1_0_30, p_1_42_43, g_1_0_18, g_2_4_7, g_0_44_44, p_0_32_32, g_1_0_4, g_1_2_3, p_0_12_12, g_2_0_25, g_0_55_55, p_0_1_1, p_0_43_43, p_0_53_53, g_0_33_33, p_0_59_59, p_0_57_57, p_1_4_5, g_4_0_55, p_2_20_23, g_2_0_9, p_2_44_47, g_0_48_48, g_5_0_31, g_0_13_13, p_0_39_39, p_1_26_27, g_1_0_48, g_2_0_37, g_0_27_27, p_0_23_23, g_0_12_12, g_3_0_27, g_0_45_45, g_1_24_25, g_6_0_63, g_1_46_47, p_0_56_56, p_1_54_55, g_1_0_40, g_1_0_28, g_1_14_15, p_1_36_37, g_0_53_53, g_3_32_39, p_0_50_50, p_1_20_21, g_2_24_27, g_1_0_60, g_1_0_14, g_0_4_4, g_0_36_36, g_2_0_21, g_0_49_49, p_1_30_31, g_1_52_53, g_1_0_2, g_4_0_39, g_3_8_15, p_0_54_54, g_0_31_31, p_0_33_33, g_2_20_23, g_5_0_47, p_0_11_11, g_4_16_31, p_2_32_35, g_2_0_33, g_1_62_63, p_0_34_34, g_2_0_57, g_0_5_5, p_0_45_45, p_1_10_11, g_1_16_17, p_0_24_24, p_3_40_47, g_1_20_21, p_0_16_16, g_1_0_24, g_0_62_62, p_1_48_49, g_3_0_43, p_2_4_7, p_0_20_20, g_0_18_18, g_0_39_39;
BlackCell U100 (.PIK(p_1_22_23), .GIK(g_1_22_23), .GKJ(g_1_20_21), .PKJ(p_1_20_21),  .GIJ(g_2_20_23), .PIJ(p_2_20_23));
BlackCell U101 (.PIK(p_1_26_27), .GIK(g_1_26_27), .GKJ(g_1_24_25), .PKJ(p_1_24_25),  .GIJ(g_2_24_27), .PIJ(p_2_24_27));
BlackCell U102 (.PIK(p_1_30_31), .GIK(g_1_30_31), .GKJ(g_1_28_29), .PKJ(p_1_28_29),  .GIJ(g_2_28_31), .PIJ(p_2_28_31));
BlackCell U103 (.PIK(p_1_34_35), .GIK(g_1_34_35), .GKJ(g_1_32_33), .PKJ(p_1_32_33),  .GIJ(g_2_32_35), .PIJ(p_2_32_35));
BlackCell U104 (.PIK(p_1_38_39), .GIK(g_1_38_39), .GKJ(g_1_36_37), .PKJ(p_1_36_37),  .GIJ(g_2_36_39), .PIJ(p_2_36_39));
BlackCell U105 (.PIK(p_1_42_43), .GIK(g_1_42_43), .GKJ(g_1_40_41), .PKJ(p_1_40_41),  .GIJ(g_2_40_43), .PIJ(p_2_40_43));
BlackCell U106 (.PIK(p_1_46_47), .GIK(g_1_46_47), .GKJ(g_1_44_45), .PKJ(p_1_44_45),  .GIJ(g_2_44_47), .PIJ(p_2_44_47));
BlackCell U107 (.PIK(p_1_50_51), .GIK(g_1_50_51), .GKJ(g_1_48_49), .PKJ(p_1_48_49),  .GIJ(g_2_48_51), .PIJ(p_2_48_51));
BlackCell U108 (.PIK(p_1_54_55), .GIK(g_1_54_55), .GKJ(g_1_52_53), .PKJ(p_1_52_53),  .GIJ(g_2_52_55), .PIJ(p_2_52_55));
BlackCell U109 (.PIK(p_1_58_59), .GIK(g_1_58_59), .GKJ(g_1_56_57), .PKJ(p_1_56_57),  .GIJ(g_2_56_59), .PIJ(p_2_56_59));
BlackCell U110 (.PIK(p_1_62_63), .GIK(g_1_62_63), .GKJ(g_1_60_61), .PKJ(p_1_60_61),  .GIJ(g_2_60_63), .PIJ(p_2_60_63));
BlackCell U112 (.PIK(p_2_12_15), .GIK(g_2_12_15), .GKJ(g_2_8_11), .PKJ(p_2_8_11),  .GIJ(g_3_8_15), .PIJ(p_3_8_15));
BlackCell U113 (.PIK(p_2_20_23), .GIK(g_2_20_23), .GKJ(g_2_16_19), .PKJ(p_2_16_19),  .GIJ(g_3_16_23), .PIJ(p_3_16_23));
BlackCell U114 (.PIK(p_2_28_31), .GIK(g_2_28_31), .GKJ(g_2_24_27), .PKJ(p_2_24_27),  .GIJ(g_3_24_31), .PIJ(p_3_24_31));
BlackCell U115 (.PIK(p_2_36_39), .GIK(g_2_36_39), .GKJ(g_2_32_35), .PKJ(p_2_32_35),  .GIJ(g_3_32_39), .PIJ(p_3_32_39));
BlackCell U116 (.PIK(p_2_44_47), .GIK(g_2_44_47), .GKJ(g_2_40_43), .PKJ(p_2_40_43),  .GIJ(g_3_40_47), .PIJ(p_3_40_47));
BlackCell U117 (.PIK(p_2_52_55), .GIK(g_2_52_55), .GKJ(g_2_48_51), .PKJ(p_2_48_51),  .GIJ(g_3_48_55), .PIJ(p_3_48_55));
BlackCell U118 (.PIK(p_2_60_63), .GIK(g_2_60_63), .GKJ(g_2_56_59), .PKJ(p_2_56_59),  .GIJ(g_3_56_63), .PIJ(p_3_56_63));
BlackCell U120 (.PIK(p_3_24_31), .GIK(g_3_24_31), .GKJ(g_3_16_23), .PKJ(p_3_16_23),  .GIJ(g_4_16_31), .PIJ(p_4_16_31));
BlackCell U121 (.PIK(p_3_40_47), .GIK(g_3_40_47), .GKJ(g_3_32_39), .PKJ(p_3_32_39),  .GIJ(g_4_32_47), .PIJ(p_4_32_47));
BlackCell U122 (.PIK(p_3_56_63), .GIK(g_3_56_63), .GKJ(g_3_48_55), .PKJ(p_3_48_55),  .GIJ(g_4_48_63), .PIJ(p_4_48_63));
BlackCell U124 (.PIK(p_4_48_63), .GIK(g_4_48_63), .GKJ(g_4_32_47), .PKJ(p_4_32_47),  .GIJ(g_5_32_63), .PIJ(p_5_32_63));
BlackCell U64 (.PIK(p_0_3_3), .GIK(g_0_3_3), .GKJ(g_0_2_2), .PKJ(p_0_2_2),  .GIJ(g_1_2_3), .PIJ(p_1_2_3));
BlackCell U65 (.PIK(p_0_5_5), .GIK(g_0_5_5), .GKJ(g_0_4_4), .PKJ(p_0_4_4),  .GIJ(g_1_4_5), .PIJ(p_1_4_5));
BlackCell U66 (.PIK(p_0_7_7), .GIK(g_0_7_7), .GKJ(g_0_6_6), .PKJ(p_0_6_6),  .GIJ(g_1_6_7), .PIJ(p_1_6_7));
BlackCell U67 (.PIK(p_0_9_9), .GIK(g_0_9_9), .GKJ(g_0_8_8), .PKJ(p_0_8_8),  .GIJ(g_1_8_9), .PIJ(p_1_8_9));
BlackCell U68 (.PIK(p_0_11_11), .GIK(g_0_11_11), .GKJ(g_0_10_10), .PKJ(p_0_10_10),  .GIJ(g_1_10_11), .PIJ(p_1_10_11));
BlackCell U69 (.PIK(p_0_13_13), .GIK(g_0_13_13), .GKJ(g_0_12_12), .PKJ(p_0_12_12),  .GIJ(g_1_12_13), .PIJ(p_1_12_13));
BlackCell U70 (.PIK(p_0_15_15), .GIK(g_0_15_15), .GKJ(g_0_14_14), .PKJ(p_0_14_14),  .GIJ(g_1_14_15), .PIJ(p_1_14_15));
BlackCell U71 (.PIK(p_0_17_17), .GIK(g_0_17_17), .GKJ(g_0_16_16), .PKJ(p_0_16_16),  .GIJ(g_1_16_17), .PIJ(p_1_16_17));
BlackCell U72 (.PIK(p_0_19_19), .GIK(g_0_19_19), .GKJ(g_0_18_18), .PKJ(p_0_18_18),  .GIJ(g_1_18_19), .PIJ(p_1_18_19));
BlackCell U73 (.PIK(p_0_21_21), .GIK(g_0_21_21), .GKJ(g_0_20_20), .PKJ(p_0_20_20),  .GIJ(g_1_20_21), .PIJ(p_1_20_21));
BlackCell U74 (.PIK(p_0_23_23), .GIK(g_0_23_23), .GKJ(g_0_22_22), .PKJ(p_0_22_22),  .GIJ(g_1_22_23), .PIJ(p_1_22_23));
BlackCell U75 (.PIK(p_0_25_25), .GIK(g_0_25_25), .GKJ(g_0_24_24), .PKJ(p_0_24_24),  .GIJ(g_1_24_25), .PIJ(p_1_24_25));
BlackCell U76 (.PIK(p_0_27_27), .GIK(g_0_27_27), .GKJ(g_0_26_26), .PKJ(p_0_26_26),  .GIJ(g_1_26_27), .PIJ(p_1_26_27));
BlackCell U77 (.PIK(p_0_29_29), .GIK(g_0_29_29), .GKJ(g_0_28_28), .PKJ(p_0_28_28),  .GIJ(g_1_28_29), .PIJ(p_1_28_29));
BlackCell U78 (.PIK(p_0_31_31), .GIK(g_0_31_31), .GKJ(g_0_30_30), .PKJ(p_0_30_30),  .GIJ(g_1_30_31), .PIJ(p_1_30_31));
BlackCell U79 (.PIK(p_0_33_33), .GIK(g_0_33_33), .GKJ(g_0_32_32), .PKJ(p_0_32_32),  .GIJ(g_1_32_33), .PIJ(p_1_32_33));
BlackCell U80 (.PIK(p_0_35_35), .GIK(g_0_35_35), .GKJ(g_0_34_34), .PKJ(p_0_34_34),  .GIJ(g_1_34_35), .PIJ(p_1_34_35));
BlackCell U81 (.PIK(p_0_37_37), .GIK(g_0_37_37), .GKJ(g_0_36_36), .PKJ(p_0_36_36),  .GIJ(g_1_36_37), .PIJ(p_1_36_37));
BlackCell U82 (.PIK(p_0_39_39), .GIK(g_0_39_39), .GKJ(g_0_38_38), .PKJ(p_0_38_38),  .GIJ(g_1_38_39), .PIJ(p_1_38_39));
BlackCell U83 (.PIK(p_0_41_41), .GIK(g_0_41_41), .GKJ(g_0_40_40), .PKJ(p_0_40_40),  .GIJ(g_1_40_41), .PIJ(p_1_40_41));
BlackCell U84 (.PIK(p_0_43_43), .GIK(g_0_43_43), .GKJ(g_0_42_42), .PKJ(p_0_42_42),  .GIJ(g_1_42_43), .PIJ(p_1_42_43));
BlackCell U85 (.PIK(p_0_45_45), .GIK(g_0_45_45), .GKJ(g_0_44_44), .PKJ(p_0_44_44),  .GIJ(g_1_44_45), .PIJ(p_1_44_45));
BlackCell U86 (.PIK(p_0_47_47), .GIK(g_0_47_47), .GKJ(g_0_46_46), .PKJ(p_0_46_46),  .GIJ(g_1_46_47), .PIJ(p_1_46_47));
BlackCell U87 (.PIK(p_0_49_49), .GIK(g_0_49_49), .GKJ(g_0_48_48), .PKJ(p_0_48_48),  .GIJ(g_1_48_49), .PIJ(p_1_48_49));
BlackCell U88 (.PIK(p_0_51_51), .GIK(g_0_51_51), .GKJ(g_0_50_50), .PKJ(p_0_50_50),  .GIJ(g_1_50_51), .PIJ(p_1_50_51));
BlackCell U89 (.PIK(p_0_53_53), .GIK(g_0_53_53), .GKJ(g_0_52_52), .PKJ(p_0_52_52),  .GIJ(g_1_52_53), .PIJ(p_1_52_53));
BlackCell U90 (.PIK(p_0_55_55), .GIK(g_0_55_55), .GKJ(g_0_54_54), .PKJ(p_0_54_54),  .GIJ(g_1_54_55), .PIJ(p_1_54_55));
BlackCell U91 (.PIK(p_0_57_57), .GIK(g_0_57_57), .GKJ(g_0_56_56), .PKJ(p_0_56_56),  .GIJ(g_1_56_57), .PIJ(p_1_56_57));
BlackCell U92 (.PIK(p_0_59_59), .GIK(g_0_59_59), .GKJ(g_0_58_58), .PKJ(p_0_58_58),  .GIJ(g_1_58_59), .PIJ(p_1_58_59));
BlackCell U93 (.PIK(p_0_61_61), .GIK(g_0_61_61), .GKJ(g_0_60_60), .PKJ(p_0_60_60),  .GIJ(g_1_60_61), .PIJ(p_1_60_61));
BlackCell U94 (.PIK(p_0_63_63), .GIK(g_0_63_63), .GKJ(g_0_62_62), .PKJ(p_0_62_62),  .GIJ(g_1_62_63), .PIJ(p_1_62_63));
BlackCell U96 (.PIK(p_1_6_7), .GIK(g_1_6_7), .GKJ(g_1_4_5), .PKJ(p_1_4_5),  .GIJ(g_2_4_7), .PIJ(p_2_4_7));
BlackCell U97 (.PIK(p_1_10_11), .GIK(g_1_10_11), .GKJ(g_1_8_9), .PKJ(p_1_8_9),  .GIJ(g_2_8_11), .PIJ(p_2_8_11));
BlackCell U98 (.PIK(p_1_14_15), .GIK(g_1_14_15), .GKJ(g_1_12_13), .PKJ(p_1_12_13),  .GIJ(g_2_12_15), .PIJ(p_2_12_15));
BlackCell U99 (.PIK(p_1_18_19), .GIK(g_1_18_19), .GKJ(g_1_16_17), .PKJ(p_1_16_17),  .GIJ(g_2_16_19), .PIJ(p_2_16_19));
GPCell UGP0 (.A(A[0]), .B(B[0]), .G(g_0_0_0), .P(p_0_0_0));
GPCell UGP1 (.A(A[1]), .B(B[1]), .G(g_0_1_1), .P(p_0_1_1));
GPCell UGP10 (.A(A[10]), .B(B[10]), .G(g_0_10_10), .P(p_0_10_10));
GPCell UGP11 (.A(A[11]), .B(B[11]), .G(g_0_11_11), .P(p_0_11_11));
GPCell UGP12 (.A(A[12]), .B(B[12]), .G(g_0_12_12), .P(p_0_12_12));
GPCell UGP13 (.A(A[13]), .B(B[13]), .G(g_0_13_13), .P(p_0_13_13));
GPCell UGP14 (.A(A[14]), .B(B[14]), .G(g_0_14_14), .P(p_0_14_14));
GPCell UGP15 (.A(A[15]), .B(B[15]), .G(g_0_15_15), .P(p_0_15_15));
GPCell UGP16 (.A(A[16]), .B(B[16]), .G(g_0_16_16), .P(p_0_16_16));
GPCell UGP17 (.A(A[17]), .B(B[17]), .G(g_0_17_17), .P(p_0_17_17));
GPCell UGP18 (.A(A[18]), .B(B[18]), .G(g_0_18_18), .P(p_0_18_18));
GPCell UGP19 (.A(A[19]), .B(B[19]), .G(g_0_19_19), .P(p_0_19_19));
GPCell UGP2 (.A(A[2]), .B(B[2]), .G(g_0_2_2), .P(p_0_2_2));
GPCell UGP20 (.A(A[20]), .B(B[20]), .G(g_0_20_20), .P(p_0_20_20));
GPCell UGP21 (.A(A[21]), .B(B[21]), .G(g_0_21_21), .P(p_0_21_21));
GPCell UGP22 (.A(A[22]), .B(B[22]), .G(g_0_22_22), .P(p_0_22_22));
GPCell UGP23 (.A(A[23]), .B(B[23]), .G(g_0_23_23), .P(p_0_23_23));
GPCell UGP24 (.A(A[24]), .B(B[24]), .G(g_0_24_24), .P(p_0_24_24));
GPCell UGP25 (.A(A[25]), .B(B[25]), .G(g_0_25_25), .P(p_0_25_25));
GPCell UGP26 (.A(A[26]), .B(B[26]), .G(g_0_26_26), .P(p_0_26_26));
GPCell UGP27 (.A(A[27]), .B(B[27]), .G(g_0_27_27), .P(p_0_27_27));
GPCell UGP28 (.A(A[28]), .B(B[28]), .G(g_0_28_28), .P(p_0_28_28));
GPCell UGP29 (.A(A[29]), .B(B[29]), .G(g_0_29_29), .P(p_0_29_29));
GPCell UGP3 (.A(A[3]), .B(B[3]), .G(g_0_3_3), .P(p_0_3_3));
GPCell UGP30 (.A(A[30]), .B(B[30]), .G(g_0_30_30), .P(p_0_30_30));
GPCell UGP31 (.A(A[31]), .B(B[31]), .G(g_0_31_31), .P(p_0_31_31));
GPCell UGP32 (.A(A[32]), .B(B[32]), .G(g_0_32_32), .P(p_0_32_32));
GPCell UGP33 (.A(A[33]), .B(B[33]), .G(g_0_33_33), .P(p_0_33_33));
GPCell UGP34 (.A(A[34]), .B(B[34]), .G(g_0_34_34), .P(p_0_34_34));
GPCell UGP35 (.A(A[35]), .B(B[35]), .G(g_0_35_35), .P(p_0_35_35));
GPCell UGP36 (.A(A[36]), .B(B[36]), .G(g_0_36_36), .P(p_0_36_36));
GPCell UGP37 (.A(A[37]), .B(B[37]), .G(g_0_37_37), .P(p_0_37_37));
GPCell UGP38 (.A(A[38]), .B(B[38]), .G(g_0_38_38), .P(p_0_38_38));
GPCell UGP39 (.A(A[39]), .B(B[39]), .G(g_0_39_39), .P(p_0_39_39));
GPCell UGP4 (.A(A[4]), .B(B[4]), .G(g_0_4_4), .P(p_0_4_4));
GPCell UGP40 (.A(A[40]), .B(B[40]), .G(g_0_40_40), .P(p_0_40_40));
GPCell UGP41 (.A(A[41]), .B(B[41]), .G(g_0_41_41), .P(p_0_41_41));
GPCell UGP42 (.A(A[42]), .B(B[42]), .G(g_0_42_42), .P(p_0_42_42));
GPCell UGP43 (.A(A[43]), .B(B[43]), .G(g_0_43_43), .P(p_0_43_43));
GPCell UGP44 (.A(A[44]), .B(B[44]), .G(g_0_44_44), .P(p_0_44_44));
GPCell UGP45 (.A(A[45]), .B(B[45]), .G(g_0_45_45), .P(p_0_45_45));
GPCell UGP46 (.A(A[46]), .B(B[46]), .G(g_0_46_46), .P(p_0_46_46));
GPCell UGP47 (.A(A[47]), .B(B[47]), .G(g_0_47_47), .P(p_0_47_47));
GPCell UGP48 (.A(A[48]), .B(B[48]), .G(g_0_48_48), .P(p_0_48_48));
GPCell UGP49 (.A(A[49]), .B(B[49]), .G(g_0_49_49), .P(p_0_49_49));
GPCell UGP5 (.A(A[5]), .B(B[5]), .G(g_0_5_5), .P(p_0_5_5));
GPCell UGP50 (.A(A[50]), .B(B[50]), .G(g_0_50_50), .P(p_0_50_50));
GPCell UGP51 (.A(A[51]), .B(B[51]), .G(g_0_51_51), .P(p_0_51_51));
GPCell UGP52 (.A(A[52]), .B(B[52]), .G(g_0_52_52), .P(p_0_52_52));
GPCell UGP53 (.A(A[53]), .B(B[53]), .G(g_0_53_53), .P(p_0_53_53));
GPCell UGP54 (.A(A[54]), .B(B[54]), .G(g_0_54_54), .P(p_0_54_54));
GPCell UGP55 (.A(A[55]), .B(B[55]), .G(g_0_55_55), .P(p_0_55_55));
GPCell UGP56 (.A(A[56]), .B(B[56]), .G(g_0_56_56), .P(p_0_56_56));
GPCell UGP57 (.A(A[57]), .B(B[57]), .G(g_0_57_57), .P(p_0_57_57));
GPCell UGP58 (.A(A[58]), .B(B[58]), .G(g_0_58_58), .P(p_0_58_58));
GPCell UGP59 (.A(A[59]), .B(B[59]), .G(g_0_59_59), .P(p_0_59_59));
GPCell UGP6 (.A(A[6]), .B(B[6]), .G(g_0_6_6), .P(p_0_6_6));
GPCell UGP60 (.A(A[60]), .B(B[60]), .G(g_0_60_60), .P(p_0_60_60));
GPCell UGP61 (.A(A[61]), .B(B[61]), .G(g_0_61_61), .P(p_0_61_61));
GPCell UGP62 (.A(A[62]), .B(B[62]), .G(g_0_62_62), .P(p_0_62_62));
GPCell UGP63 (.A(A[63]), .B(B[63]), .G(g_0_63_63), .P(p_0_63_63));
GPCell UGP7 (.A(A[7]), .B(B[7]), .G(g_0_7_7), .P(p_0_7_7));
GPCell UGP8 (.A(A[8]), .B(B[8]), .G(g_0_8_8), .P(p_0_8_8));
GPCell UGP9 (.A(A[9]), .B(B[9]), .G(g_0_9_9), .P(p_0_9_9));
GrayCell U111 (.PIK(p_2_4_7), .GIK(g_2_4_7), .GKJ(g_2_0_3), .GIJ(g_3_0_7));
GrayCell U119 (.PIK(p_3_8_15), .GIK(g_3_8_15), .GKJ(g_3_0_7), .GIJ(g_4_0_15));
GrayCell U123 (.PIK(p_4_16_31), .GIK(g_4_16_31), .GKJ(g_4_0_15), .GIJ(g_5_0_31));
GrayCell U125 (.PIK(p_5_32_63), .GIK(g_5_32_63), .GKJ(g_5_0_31), .GIJ(g_6_0_63));
GrayCell U126 (.PIK(p_4_32_47), .GIK(g_4_32_47), .GKJ(g_5_0_31), .GIJ(g_5_0_47));
GrayCell U127 (.PIK(p_3_16_23), .GIK(g_3_16_23), .GKJ(g_4_0_15), .GIJ(g_4_0_23));
GrayCell U128 (.PIK(p_3_32_39), .GIK(g_3_32_39), .GKJ(g_5_0_31), .GIJ(g_4_0_39));
GrayCell U129 (.PIK(p_3_48_55), .GIK(g_3_48_55), .GKJ(g_5_0_47), .GIJ(g_4_0_55));
GrayCell U130 (.PIK(p_2_8_11), .GIK(g_2_8_11), .GKJ(g_3_0_7), .GIJ(g_3_0_11));
GrayCell U131 (.PIK(p_2_16_19), .GIK(g_2_16_19), .GKJ(g_4_0_15), .GIJ(g_3_0_19));
GrayCell U132 (.PIK(p_2_24_27), .GIK(g_2_24_27), .GKJ(g_4_0_23), .GIJ(g_3_0_27));
GrayCell U133 (.PIK(p_2_32_35), .GIK(g_2_32_35), .GKJ(g_5_0_31), .GIJ(g_3_0_35));
GrayCell U134 (.PIK(p_2_40_43), .GIK(g_2_40_43), .GKJ(g_4_0_39), .GIJ(g_3_0_43));
GrayCell U135 (.PIK(p_2_48_51), .GIK(g_2_48_51), .GKJ(g_5_0_47), .GIJ(g_3_0_51));
GrayCell U136 (.PIK(p_2_56_59), .GIK(g_2_56_59), .GKJ(g_4_0_55), .GIJ(g_3_0_59));
GrayCell U137 (.PIK(p_1_4_5), .GIK(g_1_4_5), .GKJ(g_2_0_3), .GIJ(g_2_0_5));
GrayCell U138 (.PIK(p_1_8_9), .GIK(g_1_8_9), .GKJ(g_3_0_7), .GIJ(g_2_0_9));
GrayCell U139 (.PIK(p_1_12_13), .GIK(g_1_12_13), .GKJ(g_3_0_11), .GIJ(g_2_0_13));
GrayCell U140 (.PIK(p_1_16_17), .GIK(g_1_16_17), .GKJ(g_4_0_15), .GIJ(g_2_0_17));
GrayCell U141 (.PIK(p_1_20_21), .GIK(g_1_20_21), .GKJ(g_3_0_19), .GIJ(g_2_0_21));
GrayCell U142 (.PIK(p_1_24_25), .GIK(g_1_24_25), .GKJ(g_4_0_23), .GIJ(g_2_0_25));
GrayCell U143 (.PIK(p_1_28_29), .GIK(g_1_28_29), .GKJ(g_3_0_27), .GIJ(g_2_0_29));
GrayCell U144 (.PIK(p_1_32_33), .GIK(g_1_32_33), .GKJ(g_5_0_31), .GIJ(g_2_0_33));
GrayCell U145 (.PIK(p_1_36_37), .GIK(g_1_36_37), .GKJ(g_3_0_35), .GIJ(g_2_0_37));
GrayCell U146 (.PIK(p_1_40_41), .GIK(g_1_40_41), .GKJ(g_4_0_39), .GIJ(g_2_0_41));
GrayCell U147 (.PIK(p_1_44_45), .GIK(g_1_44_45), .GKJ(g_3_0_43), .GIJ(g_2_0_45));
GrayCell U148 (.PIK(p_1_48_49), .GIK(g_1_48_49), .GKJ(g_5_0_47), .GIJ(g_2_0_49));
GrayCell U149 (.PIK(p_1_52_53), .GIK(g_1_52_53), .GKJ(g_3_0_51), .GIJ(g_2_0_53));
GrayCell U150 (.PIK(p_1_56_57), .GIK(g_1_56_57), .GKJ(g_4_0_55), .GIJ(g_2_0_57));
GrayCell U151 (.PIK(p_1_60_61), .GIK(g_1_60_61), .GKJ(g_3_0_59), .GIJ(g_2_0_61));
GrayCell U152 (.PIK(p_0_2_2), .GIK(g_0_2_2), .GKJ(g_1_0_1), .GIJ(g_1_0_2));
GrayCell U153 (.PIK(p_0_4_4), .GIK(g_0_4_4), .GKJ(g_2_0_3), .GIJ(g_1_0_4));
GrayCell U154 (.PIK(p_0_6_6), .GIK(g_0_6_6), .GKJ(g_2_0_5), .GIJ(g_1_0_6));
GrayCell U155 (.PIK(p_0_8_8), .GIK(g_0_8_8), .GKJ(g_3_0_7), .GIJ(g_1_0_8));
GrayCell U156 (.PIK(p_0_10_10), .GIK(g_0_10_10), .GKJ(g_2_0_9), .GIJ(g_1_0_10));
GrayCell U157 (.PIK(p_0_12_12), .GIK(g_0_12_12), .GKJ(g_3_0_11), .GIJ(g_1_0_12));
GrayCell U158 (.PIK(p_0_14_14), .GIK(g_0_14_14), .GKJ(g_2_0_13), .GIJ(g_1_0_14));
GrayCell U159 (.PIK(p_0_16_16), .GIK(g_0_16_16), .GKJ(g_4_0_15), .GIJ(g_1_0_16));
GrayCell U160 (.PIK(p_0_18_18), .GIK(g_0_18_18), .GKJ(g_2_0_17), .GIJ(g_1_0_18));
GrayCell U161 (.PIK(p_0_20_20), .GIK(g_0_20_20), .GKJ(g_3_0_19), .GIJ(g_1_0_20));
GrayCell U162 (.PIK(p_0_22_22), .GIK(g_0_22_22), .GKJ(g_2_0_21), .GIJ(g_1_0_22));
GrayCell U163 (.PIK(p_0_24_24), .GIK(g_0_24_24), .GKJ(g_4_0_23), .GIJ(g_1_0_24));
GrayCell U164 (.PIK(p_0_26_26), .GIK(g_0_26_26), .GKJ(g_2_0_25), .GIJ(g_1_0_26));
GrayCell U165 (.PIK(p_0_28_28), .GIK(g_0_28_28), .GKJ(g_3_0_27), .GIJ(g_1_0_28));
GrayCell U166 (.PIK(p_0_30_30), .GIK(g_0_30_30), .GKJ(g_2_0_29), .GIJ(g_1_0_30));
GrayCell U167 (.PIK(p_0_32_32), .GIK(g_0_32_32), .GKJ(g_5_0_31), .GIJ(g_1_0_32));
GrayCell U168 (.PIK(p_0_34_34), .GIK(g_0_34_34), .GKJ(g_2_0_33), .GIJ(g_1_0_34));
GrayCell U169 (.PIK(p_0_36_36), .GIK(g_0_36_36), .GKJ(g_3_0_35), .GIJ(g_1_0_36));
GrayCell U170 (.PIK(p_0_38_38), .GIK(g_0_38_38), .GKJ(g_2_0_37), .GIJ(g_1_0_38));
GrayCell U171 (.PIK(p_0_40_40), .GIK(g_0_40_40), .GKJ(g_4_0_39), .GIJ(g_1_0_40));
GrayCell U172 (.PIK(p_0_42_42), .GIK(g_0_42_42), .GKJ(g_2_0_41), .GIJ(g_1_0_42));
GrayCell U173 (.PIK(p_0_44_44), .GIK(g_0_44_44), .GKJ(g_3_0_43), .GIJ(g_1_0_44));
GrayCell U174 (.PIK(p_0_46_46), .GIK(g_0_46_46), .GKJ(g_2_0_45), .GIJ(g_1_0_46));
GrayCell U175 (.PIK(p_0_48_48), .GIK(g_0_48_48), .GKJ(g_5_0_47), .GIJ(g_1_0_48));
GrayCell U176 (.PIK(p_0_50_50), .GIK(g_0_50_50), .GKJ(g_2_0_49), .GIJ(g_1_0_50));
GrayCell U177 (.PIK(p_0_52_52), .GIK(g_0_52_52), .GKJ(g_3_0_51), .GIJ(g_1_0_52));
GrayCell U178 (.PIK(p_0_54_54), .GIK(g_0_54_54), .GKJ(g_2_0_53), .GIJ(g_1_0_54));
GrayCell U179 (.PIK(p_0_56_56), .GIK(g_0_56_56), .GKJ(g_4_0_55), .GIJ(g_1_0_56));
GrayCell U180 (.PIK(p_0_58_58), .GIK(g_0_58_58), .GKJ(g_2_0_57), .GIJ(g_1_0_58));
GrayCell U181 (.PIK(p_0_60_60), .GIK(g_0_60_60), .GKJ(g_3_0_59), .GIJ(g_1_0_60));
GrayCell U182 (.PIK(p_0_62_62), .GIK(g_0_62_62), .GKJ(g_2_0_61), .GIJ(g_1_0_62));
GrayCell U63 (.PIK(p_0_1_1), .GIK(g_0_1_1), .GKJ(g_0_0_0), .GIJ(g_1_0_1));
GrayCell U95 (.PIK(p_1_2_3), .GIK(g_1_2_3), .GKJ(g_1_0_1), .GIJ(g_2_0_3));
assign S[64] = c[64];
assign c[0] = 1'b0;
assign c[10] = g_2_0_9;
assign c[11] = g_1_0_10;
assign c[12] = g_3_0_11;
assign c[13] = g_1_0_12;
assign c[14] = g_2_0_13;
assign c[15] = g_1_0_14;
assign c[16] = g_4_0_15;
assign c[17] = g_1_0_16;
assign c[18] = g_2_0_17;
assign c[19] = g_1_0_18;
assign c[1] = g_0_0_0;
assign c[20] = g_3_0_19;
assign c[21] = g_1_0_20;
assign c[22] = g_2_0_21;
assign c[23] = g_1_0_22;
assign c[24] = g_4_0_23;
assign c[25] = g_1_0_24;
assign c[26] = g_2_0_25;
assign c[27] = g_1_0_26;
assign c[28] = g_3_0_27;
assign c[29] = g_1_0_28;
assign c[2] = g_1_0_1;
assign c[30] = g_2_0_29;
assign c[31] = g_1_0_30;
assign c[32] = g_5_0_31;
assign c[33] = g_1_0_32;
assign c[34] = g_2_0_33;
assign c[35] = g_1_0_34;
assign c[36] = g_3_0_35;
assign c[37] = g_1_0_36;
assign c[38] = g_2_0_37;
assign c[39] = g_1_0_38;
assign c[3] = g_1_0_2;
assign c[40] = g_4_0_39;
assign c[41] = g_1_0_40;
assign c[42] = g_2_0_41;
assign c[43] = g_1_0_42;
assign c[44] = g_3_0_43;
assign c[45] = g_1_0_44;
assign c[46] = g_2_0_45;
assign c[47] = g_1_0_46;
assign c[48] = g_5_0_47;
assign c[49] = g_1_0_48;
assign c[4] = g_2_0_3;
assign c[50] = g_2_0_49;
assign c[51] = g_1_0_50;
assign c[52] = g_3_0_51;
assign c[53] = g_1_0_52;
assign c[54] = g_2_0_53;
assign c[55] = g_1_0_54;
assign c[56] = g_4_0_55;
assign c[57] = g_1_0_56;
assign c[58] = g_2_0_57;
assign c[59] = g_1_0_58;
assign c[5] = g_1_0_4;
assign c[60] = g_3_0_59;
assign c[61] = g_1_0_60;
assign c[62] = g_2_0_61;
assign c[63] = g_1_0_62;
assign c[64] = g_6_0_63;
assign c[6] = g_2_0_5;
assign c[7] = g_1_0_6;
assign c[8] = g_3_0_7;
assign c[9] = g_1_0_8;
xor UXOR0 (S[0], p_0_0_0, c[0]);
xor UXOR1 (S[1], p_0_1_1, c[1]);
xor UXOR10 (S[10], p_0_10_10, c[10]);
xor UXOR11 (S[11], p_0_11_11, c[11]);
xor UXOR12 (S[12], p_0_12_12, c[12]);
xor UXOR13 (S[13], p_0_13_13, c[13]);
xor UXOR14 (S[14], p_0_14_14, c[14]);
xor UXOR15 (S[15], p_0_15_15, c[15]);
xor UXOR16 (S[16], p_0_16_16, c[16]);
xor UXOR17 (S[17], p_0_17_17, c[17]);
xor UXOR18 (S[18], p_0_18_18, c[18]);
xor UXOR19 (S[19], p_0_19_19, c[19]);
xor UXOR2 (S[2], p_0_2_2, c[2]);
xor UXOR20 (S[20], p_0_20_20, c[20]);
xor UXOR21 (S[21], p_0_21_21, c[21]);
xor UXOR22 (S[22], p_0_22_22, c[22]);
xor UXOR23 (S[23], p_0_23_23, c[23]);
xor UXOR24 (S[24], p_0_24_24, c[24]);
xor UXOR25 (S[25], p_0_25_25, c[25]);
xor UXOR26 (S[26], p_0_26_26, c[26]);
xor UXOR27 (S[27], p_0_27_27, c[27]);
xor UXOR28 (S[28], p_0_28_28, c[28]);
xor UXOR29 (S[29], p_0_29_29, c[29]);
xor UXOR3 (S[3], p_0_3_3, c[3]);
xor UXOR30 (S[30], p_0_30_30, c[30]);
xor UXOR31 (S[31], p_0_31_31, c[31]);
xor UXOR32 (S[32], p_0_32_32, c[32]);
xor UXOR33 (S[33], p_0_33_33, c[33]);
xor UXOR34 (S[34], p_0_34_34, c[34]);
xor UXOR35 (S[35], p_0_35_35, c[35]);
xor UXOR36 (S[36], p_0_36_36, c[36]);
xor UXOR37 (S[37], p_0_37_37, c[37]);
xor UXOR38 (S[38], p_0_38_38, c[38]);
xor UXOR39 (S[39], p_0_39_39, c[39]);
xor UXOR4 (S[4], p_0_4_4, c[4]);
xor UXOR40 (S[40], p_0_40_40, c[40]);
xor UXOR41 (S[41], p_0_41_41, c[41]);
xor UXOR42 (S[42], p_0_42_42, c[42]);
xor UXOR43 (S[43], p_0_43_43, c[43]);
xor UXOR44 (S[44], p_0_44_44, c[44]);
xor UXOR45 (S[45], p_0_45_45, c[45]);
xor UXOR46 (S[46], p_0_46_46, c[46]);
xor UXOR47 (S[47], p_0_47_47, c[47]);
xor UXOR48 (S[48], p_0_48_48, c[48]);
xor UXOR49 (S[49], p_0_49_49, c[49]);
xor UXOR5 (S[5], p_0_5_5, c[5]);
xor UXOR50 (S[50], p_0_50_50, c[50]);
xor UXOR51 (S[51], p_0_51_51, c[51]);
xor UXOR52 (S[52], p_0_52_52, c[52]);
xor UXOR53 (S[53], p_0_53_53, c[53]);
xor UXOR54 (S[54], p_0_54_54, c[54]);
xor UXOR55 (S[55], p_0_55_55, c[55]);
xor UXOR56 (S[56], p_0_56_56, c[56]);
xor UXOR57 (S[57], p_0_57_57, c[57]);
xor UXOR58 (S[58], p_0_58_58, c[58]);
xor UXOR59 (S[59], p_0_59_59, c[59]);
xor UXOR6 (S[6], p_0_6_6, c[6]);
xor UXOR60 (S[60], p_0_60_60, c[60]);
xor UXOR61 (S[61], p_0_61_61, c[61]);
xor UXOR62 (S[62], p_0_62_62, c[62]);
xor UXOR63 (S[63], p_0_63_63, c[63]);
xor UXOR7 (S[7], p_0_7_7, c[7]);
xor UXOR8 (S[8], p_0_8_8, c[8]);
xor UXOR9 (S[9], p_0_9_9, c[9]);
endmodule