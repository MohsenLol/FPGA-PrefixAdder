library verilog;
use verilog.vl_types.all;
entity rippleCarry2b_tb is
end rippleCarry2b_tb;
