`timescale 1ns/1ns
module testbench;
wire [_N_ : 0] S;
reg [_N_ - 1 : 0] A, B;
reg [_N_ : 0] SR;
_X_ UUT(.A(A), .B(B), .S(S));
reg condi, condj;
integer errors = 0;
initial begin
    condi = 1;
    condj = 1;
    A = _S_;
    B = _S_;
    while(condi) begin
        condj = 1;
        while(condj) begin
            SR = A + B;
            #1;
            if(S !== SR) begin
                errors = errors + 1;
                $display("Missmatch : %dD(%bB) + %dD(%bB) => %dD(%bB) != %dD", A, A, B, B, S, S, SR);
            end 
            B = B + 1;
            if(B == _E_) begin
                condj = 0;
            end
        end
        A = A + 1;
        if(A == _E_) begin 
            condi = 0;
        end

    end
    $display("Total Error count is %d", errors);
    $stop();
end
endmodule