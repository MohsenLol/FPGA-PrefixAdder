library verilog;
use verilog.vl_types.all;
entity BrentKung8b_tb is
end BrentKung8b_tb;
