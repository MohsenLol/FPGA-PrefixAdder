library verilog;
use verilog.vl_types.all;
entity LadnerFischer8b_tb is
end LadnerFischer8b_tb;
