library verilog;
use verilog.vl_types.all;
entity BrentKung32b_etb is
end BrentKung32b_etb;
