module BrentKung32b (A, B, S);
input [31 : 0] A;
input [31 : 0] B;
output [32 : 0] S;
wire p_1_4_5, p_1_8_9, g_2_0_29, p_0_14_14, g_2_28_31, g_2_16_19, p_4_16_31, c [32 : 0], g_0_20_20, p_2_20_23, g_0_25_25, g_2_0_9, p_0_26_26, g_3_0_11, p_2_12_15, p_0_18_18, g_5_0_31, p_1_14_15, g_0_13_13, g_0_8_8, p_1_26_27, g_1_12_13, p_3_24_31, p_0_4_4, g_0_21_21, g_1_0_22, g_1_0_8, g_0_27_27, p_0_23_23, g_0_12_12, g_0_2_2, g_1_28_29, p_2_16_19, p_0_15_15, g_3_0_27, p_0_31_31, g_1_24_25, g_3_24_31, g_4_0_15, g_0_19_19, p_1_12_13, g_2_0_13, g_0_22_22, p_2_28_31, g_0_11_11, g_0_23_23, p_0_13_13, p_2_24_27, p_1_16_17, p_0_25_25, p_0_9_9, g_2_0_3, g_1_0_28, g_1_14_15, g_0_17_17, p_0_29_29, g_1_0_12, p_0_21_21, g_0_30_30, g_3_0_19, p_1_20_21, g_0_15_15, p_1_28_29, g_2_24_27, p_1_24_25, g_1_0_14, g_1_0_26, g_1_6_7, g_1_0_20, g_1_0_1, g_0_4_4, g_3_16_23, g_4_0_23, p_0_8_8, p_3_16_23, p_1_18_19, g_0_9_9, g_2_0_21, p_1_30_31, g_1_0_2, p_0_3_3, p_3_8_15, g_3_8_15, p_1_6_7, g_1_10_11, g_1_22_23, p_0_19_19, p_0_6_6, p_0_17_17, p_0_0_0, g_2_8_11, p_0_2_2, g_0_31_31, g_2_20_23, p_0_11_11, p_0_10_10, g_0_29_29, g_0_7_7, g_4_16_31, g_1_18_19, g_1_4_5, p_0_7_7, g_3_0_7, g_0_6_6, g_0_10_10, g_0_0_0, g_0_3_3, g_1_26_27, g_1_0_6, g_0_26_26, g_0_1_1, p_0_22_22, g_2_0_17, g_1_8_9, p_1_22_23, p_2_8_11, g_0_28_28, g_2_0_5, g_0_5_5, p_1_10_11, p_0_30_30, g_0_24_24, g_1_16_17, p_0_24_24, g_1_0_16, g_0_16_16, g_1_20_21, g_1_30_31, p_0_27_27, g_0_14_14, g_1_0_10, p_0_16_16, p_0_5_5, g_2_12_15, g_1_0_30, g_1_0_18, g_1_0_24, g_2_4_7, p_0_28_28, p_1_2_3, g_1_0_4, g_1_2_3, p_0_12_12, p_0_20_20, p_2_4_7, g_2_0_25, g_0_18_18, p_0_1_1;
BlackCell U32 (.PIK(p_0_3_3), .GIK(g_0_3_3), .GKJ(g_0_2_2), .PKJ(p_0_2_2),  .GIJ(g_1_2_3), .PIJ(p_1_2_3));
BlackCell U33 (.PIK(p_0_5_5), .GIK(g_0_5_5), .GKJ(g_0_4_4), .PKJ(p_0_4_4),  .GIJ(g_1_4_5), .PIJ(p_1_4_5));
BlackCell U34 (.PIK(p_0_7_7), .GIK(g_0_7_7), .GKJ(g_0_6_6), .PKJ(p_0_6_6),  .GIJ(g_1_6_7), .PIJ(p_1_6_7));
BlackCell U35 (.PIK(p_0_9_9), .GIK(g_0_9_9), .GKJ(g_0_8_8), .PKJ(p_0_8_8),  .GIJ(g_1_8_9), .PIJ(p_1_8_9));
BlackCell U36 (.PIK(p_0_11_11), .GIK(g_0_11_11), .GKJ(g_0_10_10), .PKJ(p_0_10_10),  .GIJ(g_1_10_11), .PIJ(p_1_10_11));
BlackCell U37 (.PIK(p_0_13_13), .GIK(g_0_13_13), .GKJ(g_0_12_12), .PKJ(p_0_12_12),  .GIJ(g_1_12_13), .PIJ(p_1_12_13));
BlackCell U38 (.PIK(p_0_15_15), .GIK(g_0_15_15), .GKJ(g_0_14_14), .PKJ(p_0_14_14),  .GIJ(g_1_14_15), .PIJ(p_1_14_15));
BlackCell U39 (.PIK(p_0_17_17), .GIK(g_0_17_17), .GKJ(g_0_16_16), .PKJ(p_0_16_16),  .GIJ(g_1_16_17), .PIJ(p_1_16_17));
BlackCell U40 (.PIK(p_0_19_19), .GIK(g_0_19_19), .GKJ(g_0_18_18), .PKJ(p_0_18_18),  .GIJ(g_1_18_19), .PIJ(p_1_18_19));
BlackCell U41 (.PIK(p_0_21_21), .GIK(g_0_21_21), .GKJ(g_0_20_20), .PKJ(p_0_20_20),  .GIJ(g_1_20_21), .PIJ(p_1_20_21));
BlackCell U42 (.PIK(p_0_23_23), .GIK(g_0_23_23), .GKJ(g_0_22_22), .PKJ(p_0_22_22),  .GIJ(g_1_22_23), .PIJ(p_1_22_23));
BlackCell U43 (.PIK(p_0_25_25), .GIK(g_0_25_25), .GKJ(g_0_24_24), .PKJ(p_0_24_24),  .GIJ(g_1_24_25), .PIJ(p_1_24_25));
BlackCell U44 (.PIK(p_0_27_27), .GIK(g_0_27_27), .GKJ(g_0_26_26), .PKJ(p_0_26_26),  .GIJ(g_1_26_27), .PIJ(p_1_26_27));
BlackCell U45 (.PIK(p_0_29_29), .GIK(g_0_29_29), .GKJ(g_0_28_28), .PKJ(p_0_28_28),  .GIJ(g_1_28_29), .PIJ(p_1_28_29));
BlackCell U46 (.PIK(p_0_31_31), .GIK(g_0_31_31), .GKJ(g_0_30_30), .PKJ(p_0_30_30),  .GIJ(g_1_30_31), .PIJ(p_1_30_31));
BlackCell U48 (.PIK(p_1_6_7), .GIK(g_1_6_7), .GKJ(g_1_4_5), .PKJ(p_1_4_5),  .GIJ(g_2_4_7), .PIJ(p_2_4_7));
BlackCell U49 (.PIK(p_1_10_11), .GIK(g_1_10_11), .GKJ(g_1_8_9), .PKJ(p_1_8_9),  .GIJ(g_2_8_11), .PIJ(p_2_8_11));
BlackCell U50 (.PIK(p_1_14_15), .GIK(g_1_14_15), .GKJ(g_1_12_13), .PKJ(p_1_12_13),  .GIJ(g_2_12_15), .PIJ(p_2_12_15));
BlackCell U51 (.PIK(p_1_18_19), .GIK(g_1_18_19), .GKJ(g_1_16_17), .PKJ(p_1_16_17),  .GIJ(g_2_16_19), .PIJ(p_2_16_19));
BlackCell U52 (.PIK(p_1_22_23), .GIK(g_1_22_23), .GKJ(g_1_20_21), .PKJ(p_1_20_21),  .GIJ(g_2_20_23), .PIJ(p_2_20_23));
BlackCell U53 (.PIK(p_1_26_27), .GIK(g_1_26_27), .GKJ(g_1_24_25), .PKJ(p_1_24_25),  .GIJ(g_2_24_27), .PIJ(p_2_24_27));
BlackCell U54 (.PIK(p_1_30_31), .GIK(g_1_30_31), .GKJ(g_1_28_29), .PKJ(p_1_28_29),  .GIJ(g_2_28_31), .PIJ(p_2_28_31));
BlackCell U56 (.PIK(p_2_12_15), .GIK(g_2_12_15), .GKJ(g_2_8_11), .PKJ(p_2_8_11),  .GIJ(g_3_8_15), .PIJ(p_3_8_15));
BlackCell U57 (.PIK(p_2_20_23), .GIK(g_2_20_23), .GKJ(g_2_16_19), .PKJ(p_2_16_19),  .GIJ(g_3_16_23), .PIJ(p_3_16_23));
BlackCell U58 (.PIK(p_2_28_31), .GIK(g_2_28_31), .GKJ(g_2_24_27), .PKJ(p_2_24_27),  .GIJ(g_3_24_31), .PIJ(p_3_24_31));
BlackCell U60 (.PIK(p_3_24_31), .GIK(g_3_24_31), .GKJ(g_3_16_23), .PKJ(p_3_16_23),  .GIJ(g_4_16_31), .PIJ(p_4_16_31));
GPCell UGP0 (.A(A[0]), .B(B[0]), .G(g_0_0_0), .P(p_0_0_0));
GPCell UGP1 (.A(A[1]), .B(B[1]), .G(g_0_1_1), .P(p_0_1_1));
GPCell UGP10 (.A(A[10]), .B(B[10]), .G(g_0_10_10), .P(p_0_10_10));
GPCell UGP11 (.A(A[11]), .B(B[11]), .G(g_0_11_11), .P(p_0_11_11));
GPCell UGP12 (.A(A[12]), .B(B[12]), .G(g_0_12_12), .P(p_0_12_12));
GPCell UGP13 (.A(A[13]), .B(B[13]), .G(g_0_13_13), .P(p_0_13_13));
GPCell UGP14 (.A(A[14]), .B(B[14]), .G(g_0_14_14), .P(p_0_14_14));
GPCell UGP15 (.A(A[15]), .B(B[15]), .G(g_0_15_15), .P(p_0_15_15));
GPCell UGP16 (.A(A[16]), .B(B[16]), .G(g_0_16_16), .P(p_0_16_16));
GPCell UGP17 (.A(A[17]), .B(B[17]), .G(g_0_17_17), .P(p_0_17_17));
GPCell UGP18 (.A(A[18]), .B(B[18]), .G(g_0_18_18), .P(p_0_18_18));
GPCell UGP19 (.A(A[19]), .B(B[19]), .G(g_0_19_19), .P(p_0_19_19));
GPCell UGP2 (.A(A[2]), .B(B[2]), .G(g_0_2_2), .P(p_0_2_2));
GPCell UGP20 (.A(A[20]), .B(B[20]), .G(g_0_20_20), .P(p_0_20_20));
GPCell UGP21 (.A(A[21]), .B(B[21]), .G(g_0_21_21), .P(p_0_21_21));
GPCell UGP22 (.A(A[22]), .B(B[22]), .G(g_0_22_22), .P(p_0_22_22));
GPCell UGP23 (.A(A[23]), .B(B[23]), .G(g_0_23_23), .P(p_0_23_23));
GPCell UGP24 (.A(A[24]), .B(B[24]), .G(g_0_24_24), .P(p_0_24_24));
GPCell UGP25 (.A(A[25]), .B(B[25]), .G(g_0_25_25), .P(p_0_25_25));
GPCell UGP26 (.A(A[26]), .B(B[26]), .G(g_0_26_26), .P(p_0_26_26));
GPCell UGP27 (.A(A[27]), .B(B[27]), .G(g_0_27_27), .P(p_0_27_27));
GPCell UGP28 (.A(A[28]), .B(B[28]), .G(g_0_28_28), .P(p_0_28_28));
GPCell UGP29 (.A(A[29]), .B(B[29]), .G(g_0_29_29), .P(p_0_29_29));
GPCell UGP3 (.A(A[3]), .B(B[3]), .G(g_0_3_3), .P(p_0_3_3));
GPCell UGP30 (.A(A[30]), .B(B[30]), .G(g_0_30_30), .P(p_0_30_30));
GPCell UGP31 (.A(A[31]), .B(B[31]), .G(g_0_31_31), .P(p_0_31_31));
GPCell UGP4 (.A(A[4]), .B(B[4]), .G(g_0_4_4), .P(p_0_4_4));
GPCell UGP5 (.A(A[5]), .B(B[5]), .G(g_0_5_5), .P(p_0_5_5));
GPCell UGP6 (.A(A[6]), .B(B[6]), .G(g_0_6_6), .P(p_0_6_6));
GPCell UGP7 (.A(A[7]), .B(B[7]), .G(g_0_7_7), .P(p_0_7_7));
GPCell UGP8 (.A(A[8]), .B(B[8]), .G(g_0_8_8), .P(p_0_8_8));
GPCell UGP9 (.A(A[9]), .B(B[9]), .G(g_0_9_9), .P(p_0_9_9));
GrayCell U31 (.PIK(p_0_1_1), .GIK(g_0_1_1), .GKJ(g_0_0_0), .GIJ(g_1_0_1));
GrayCell U47 (.PIK(p_1_2_3), .GIK(g_1_2_3), .GKJ(g_1_0_1), .GIJ(g_2_0_3));
GrayCell U55 (.PIK(p_2_4_7), .GIK(g_2_4_7), .GKJ(g_2_0_3), .GIJ(g_3_0_7));
GrayCell U59 (.PIK(p_3_8_15), .GIK(g_3_8_15), .GKJ(g_3_0_7), .GIJ(g_4_0_15));
GrayCell U61 (.PIK(p_4_16_31), .GIK(g_4_16_31), .GKJ(g_4_0_15), .GIJ(g_5_0_31));
GrayCell U62 (.PIK(p_3_16_23), .GIK(g_3_16_23), .GKJ(g_4_0_15), .GIJ(g_4_0_23));
GrayCell U63 (.PIK(p_2_8_11), .GIK(g_2_8_11), .GKJ(g_3_0_7), .GIJ(g_3_0_11));
GrayCell U64 (.PIK(p_2_16_19), .GIK(g_2_16_19), .GKJ(g_4_0_15), .GIJ(g_3_0_19));
GrayCell U65 (.PIK(p_2_24_27), .GIK(g_2_24_27), .GKJ(g_4_0_23), .GIJ(g_3_0_27));
GrayCell U66 (.PIK(p_1_4_5), .GIK(g_1_4_5), .GKJ(g_2_0_3), .GIJ(g_2_0_5));
GrayCell U67 (.PIK(p_1_8_9), .GIK(g_1_8_9), .GKJ(g_3_0_7), .GIJ(g_2_0_9));
GrayCell U68 (.PIK(p_1_12_13), .GIK(g_1_12_13), .GKJ(g_3_0_11), .GIJ(g_2_0_13));
GrayCell U69 (.PIK(p_1_16_17), .GIK(g_1_16_17), .GKJ(g_4_0_15), .GIJ(g_2_0_17));
GrayCell U70 (.PIK(p_1_20_21), .GIK(g_1_20_21), .GKJ(g_3_0_19), .GIJ(g_2_0_21));
GrayCell U71 (.PIK(p_1_24_25), .GIK(g_1_24_25), .GKJ(g_4_0_23), .GIJ(g_2_0_25));
GrayCell U72 (.PIK(p_1_28_29), .GIK(g_1_28_29), .GKJ(g_3_0_27), .GIJ(g_2_0_29));
GrayCell U73 (.PIK(p_0_2_2), .GIK(g_0_2_2), .GKJ(g_1_0_1), .GIJ(g_1_0_2));
GrayCell U74 (.PIK(p_0_4_4), .GIK(g_0_4_4), .GKJ(g_2_0_3), .GIJ(g_1_0_4));
GrayCell U75 (.PIK(p_0_6_6), .GIK(g_0_6_6), .GKJ(g_2_0_5), .GIJ(g_1_0_6));
GrayCell U76 (.PIK(p_0_8_8), .GIK(g_0_8_8), .GKJ(g_3_0_7), .GIJ(g_1_0_8));
GrayCell U77 (.PIK(p_0_10_10), .GIK(g_0_10_10), .GKJ(g_2_0_9), .GIJ(g_1_0_10));
GrayCell U78 (.PIK(p_0_12_12), .GIK(g_0_12_12), .GKJ(g_3_0_11), .GIJ(g_1_0_12));
GrayCell U79 (.PIK(p_0_14_14), .GIK(g_0_14_14), .GKJ(g_2_0_13), .GIJ(g_1_0_14));
GrayCell U80 (.PIK(p_0_16_16), .GIK(g_0_16_16), .GKJ(g_4_0_15), .GIJ(g_1_0_16));
GrayCell U81 (.PIK(p_0_18_18), .GIK(g_0_18_18), .GKJ(g_2_0_17), .GIJ(g_1_0_18));
GrayCell U82 (.PIK(p_0_20_20), .GIK(g_0_20_20), .GKJ(g_3_0_19), .GIJ(g_1_0_20));
GrayCell U83 (.PIK(p_0_22_22), .GIK(g_0_22_22), .GKJ(g_2_0_21), .GIJ(g_1_0_22));
GrayCell U84 (.PIK(p_0_24_24), .GIK(g_0_24_24), .GKJ(g_4_0_23), .GIJ(g_1_0_24));
GrayCell U85 (.PIK(p_0_26_26), .GIK(g_0_26_26), .GKJ(g_2_0_25), .GIJ(g_1_0_26));
GrayCell U86 (.PIK(p_0_28_28), .GIK(g_0_28_28), .GKJ(g_3_0_27), .GIJ(g_1_0_28));
GrayCell U87 (.PIK(p_0_30_30), .GIK(g_0_30_30), .GKJ(g_2_0_29), .GIJ(g_1_0_30));
assign S[32] = c[32];
assign c[0] = 1'b0;
assign c[10] = g_2_0_9;
assign c[11] = g_1_0_10;
assign c[12] = g_3_0_11;
assign c[13] = g_1_0_12;
assign c[14] = g_2_0_13;
assign c[15] = g_1_0_14;
assign c[16] = g_4_0_15;
assign c[17] = g_1_0_16;
assign c[18] = g_2_0_17;
assign c[19] = g_1_0_18;
assign c[1] = g_0_0_0;
assign c[20] = g_3_0_19;
assign c[21] = g_1_0_20;
assign c[22] = g_2_0_21;
assign c[23] = g_1_0_22;
assign c[24] = g_4_0_23;
assign c[25] = g_1_0_24;
assign c[26] = g_2_0_25;
assign c[27] = g_1_0_26;
assign c[28] = g_3_0_27;
assign c[29] = g_1_0_28;
assign c[2] = g_1_0_1;
assign c[30] = g_2_0_29;
assign c[31] = g_1_0_30;
assign c[32] = g_5_0_31;
assign c[3] = g_1_0_2;
assign c[4] = g_2_0_3;
assign c[5] = g_1_0_4;
assign c[6] = g_2_0_5;
assign c[7] = g_1_0_6;
assign c[8] = g_3_0_7;
assign c[9] = g_1_0_8;
xor UXOR0 (S[0], p_0_0_0, c[0]);
xor UXOR1 (S[1], p_0_1_1, c[1]);
xor UXOR10 (S[10], p_0_10_10, c[10]);
xor UXOR11 (S[11], p_0_11_11, c[11]);
xor UXOR12 (S[12], p_0_12_12, c[12]);
xor UXOR13 (S[13], p_0_13_13, c[13]);
xor UXOR14 (S[14], p_0_14_14, c[14]);
xor UXOR15 (S[15], p_0_15_15, c[15]);
xor UXOR16 (S[16], p_0_16_16, c[16]);
xor UXOR17 (S[17], p_0_17_17, c[17]);
xor UXOR18 (S[18], p_0_18_18, c[18]);
xor UXOR19 (S[19], p_0_19_19, c[19]);
xor UXOR2 (S[2], p_0_2_2, c[2]);
xor UXOR20 (S[20], p_0_20_20, c[20]);
xor UXOR21 (S[21], p_0_21_21, c[21]);
xor UXOR22 (S[22], p_0_22_22, c[22]);
xor UXOR23 (S[23], p_0_23_23, c[23]);
xor UXOR24 (S[24], p_0_24_24, c[24]);
xor UXOR25 (S[25], p_0_25_25, c[25]);
xor UXOR26 (S[26], p_0_26_26, c[26]);
xor UXOR27 (S[27], p_0_27_27, c[27]);
xor UXOR28 (S[28], p_0_28_28, c[28]);
xor UXOR29 (S[29], p_0_29_29, c[29]);
xor UXOR3 (S[3], p_0_3_3, c[3]);
xor UXOR30 (S[30], p_0_30_30, c[30]);
xor UXOR31 (S[31], p_0_31_31, c[31]);
xor UXOR4 (S[4], p_0_4_4, c[4]);
xor UXOR5 (S[5], p_0_5_5, c[5]);
xor UXOR6 (S[6], p_0_6_6, c[6]);
xor UXOR7 (S[7], p_0_7_7, c[7]);
xor UXOR8 (S[8], p_0_8_8, c[8]);
xor UXOR9 (S[9], p_0_9_9, c[9]);
endmodule