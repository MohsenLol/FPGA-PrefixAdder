library verilog;
use verilog.vl_types.all;
entity KoggeStone32b_tb is
end KoggeStone32b_tb;
