module BrentKung16b (A, B, S);
input [15 : 0] A;
input [15 : 0] B;
output [16 : 0] S;
wire p_1_4_5, p_1_8_9, p_0_14_14, c [16 : 0], g_2_0_9, g_3_0_11, p_2_12_15, p_1_14_15, g_0_13_13, g_0_8_8, g_1_12_13, p_0_4_4, g_1_0_8, g_0_12_12, g_0_2_2, p_0_15_15, g_4_0_15, p_1_12_13, g_2_0_13, g_0_11_11, p_0_13_13, g_2_0_3, p_0_9_9, g_1_14_15, g_1_0_12, g_0_15_15, g_1_0_14, g_1_6_7, g_1_0_1, g_0_4_4, p_0_8_8, g_0_9_9, g_1_0_2, p_0_3_3, p_3_8_15, g_3_8_15, p_1_6_7, g_1_10_11, p_0_6_6, p_0_0_0, g_2_8_11, p_0_2_2, p_0_11_11, p_0_10_10, g_0_7_7, g_3_0_7, g_1_4_5, p_0_7_7, g_0_6_6, g_0_10_10, g_0_0_0, g_0_3_3, g_1_0_6, g_0_1_1, g_1_8_9, p_2_8_11, g_2_0_5, g_0_5_5, p_1_10_11, g_0_14_14, g_1_0_10, p_0_5_5, g_2_12_15, g_2_4_7, p_1_2_3, g_1_0_4, g_1_2_3, p_0_12_12, p_2_4_7, p_0_1_1;
BlackCell U16 (.PIK(p_0_3_3), .GIK(g_0_3_3), .GKJ(g_0_2_2), .PKJ(p_0_2_2),  .GIJ(g_1_2_3), .PIJ(p_1_2_3));
BlackCell U17 (.PIK(p_0_5_5), .GIK(g_0_5_5), .GKJ(g_0_4_4), .PKJ(p_0_4_4),  .GIJ(g_1_4_5), .PIJ(p_1_4_5));
BlackCell U18 (.PIK(p_0_7_7), .GIK(g_0_7_7), .GKJ(g_0_6_6), .PKJ(p_0_6_6),  .GIJ(g_1_6_7), .PIJ(p_1_6_7));
BlackCell U19 (.PIK(p_0_9_9), .GIK(g_0_9_9), .GKJ(g_0_8_8), .PKJ(p_0_8_8),  .GIJ(g_1_8_9), .PIJ(p_1_8_9));
BlackCell U20 (.PIK(p_0_11_11), .GIK(g_0_11_11), .GKJ(g_0_10_10), .PKJ(p_0_10_10),  .GIJ(g_1_10_11), .PIJ(p_1_10_11));
BlackCell U21 (.PIK(p_0_13_13), .GIK(g_0_13_13), .GKJ(g_0_12_12), .PKJ(p_0_12_12),  .GIJ(g_1_12_13), .PIJ(p_1_12_13));
BlackCell U22 (.PIK(p_0_15_15), .GIK(g_0_15_15), .GKJ(g_0_14_14), .PKJ(p_0_14_14),  .GIJ(g_1_14_15), .PIJ(p_1_14_15));
BlackCell U24 (.PIK(p_1_6_7), .GIK(g_1_6_7), .GKJ(g_1_4_5), .PKJ(p_1_4_5),  .GIJ(g_2_4_7), .PIJ(p_2_4_7));
BlackCell U25 (.PIK(p_1_10_11), .GIK(g_1_10_11), .GKJ(g_1_8_9), .PKJ(p_1_8_9),  .GIJ(g_2_8_11), .PIJ(p_2_8_11));
BlackCell U26 (.PIK(p_1_14_15), .GIK(g_1_14_15), .GKJ(g_1_12_13), .PKJ(p_1_12_13),  .GIJ(g_2_12_15), .PIJ(p_2_12_15));
BlackCell U28 (.PIK(p_2_12_15), .GIK(g_2_12_15), .GKJ(g_2_8_11), .PKJ(p_2_8_11),  .GIJ(g_3_8_15), .PIJ(p_3_8_15));
GPCell UGP0 (.A(A[0]), .B(B[0]), .G(g_0_0_0), .P(p_0_0_0));
GPCell UGP1 (.A(A[1]), .B(B[1]), .G(g_0_1_1), .P(p_0_1_1));
GPCell UGP10 (.A(A[10]), .B(B[10]), .G(g_0_10_10), .P(p_0_10_10));
GPCell UGP11 (.A(A[11]), .B(B[11]), .G(g_0_11_11), .P(p_0_11_11));
GPCell UGP12 (.A(A[12]), .B(B[12]), .G(g_0_12_12), .P(p_0_12_12));
GPCell UGP13 (.A(A[13]), .B(B[13]), .G(g_0_13_13), .P(p_0_13_13));
GPCell UGP14 (.A(A[14]), .B(B[14]), .G(g_0_14_14), .P(p_0_14_14));
GPCell UGP15 (.A(A[15]), .B(B[15]), .G(g_0_15_15), .P(p_0_15_15));
GPCell UGP2 (.A(A[2]), .B(B[2]), .G(g_0_2_2), .P(p_0_2_2));
GPCell UGP3 (.A(A[3]), .B(B[3]), .G(g_0_3_3), .P(p_0_3_3));
GPCell UGP4 (.A(A[4]), .B(B[4]), .G(g_0_4_4), .P(p_0_4_4));
GPCell UGP5 (.A(A[5]), .B(B[5]), .G(g_0_5_5), .P(p_0_5_5));
GPCell UGP6 (.A(A[6]), .B(B[6]), .G(g_0_6_6), .P(p_0_6_6));
GPCell UGP7 (.A(A[7]), .B(B[7]), .G(g_0_7_7), .P(p_0_7_7));
GPCell UGP8 (.A(A[8]), .B(B[8]), .G(g_0_8_8), .P(p_0_8_8));
GPCell UGP9 (.A(A[9]), .B(B[9]), .G(g_0_9_9), .P(p_0_9_9));
GrayCell U15 (.PIK(p_0_1_1), .GIK(g_0_1_1), .GKJ(g_0_0_0), .GIJ(g_1_0_1));
GrayCell U23 (.PIK(p_1_2_3), .GIK(g_1_2_3), .GKJ(g_1_0_1), .GIJ(g_2_0_3));
GrayCell U27 (.PIK(p_2_4_7), .GIK(g_2_4_7), .GKJ(g_2_0_3), .GIJ(g_3_0_7));
GrayCell U29 (.PIK(p_3_8_15), .GIK(g_3_8_15), .GKJ(g_3_0_7), .GIJ(g_4_0_15));
GrayCell U30 (.PIK(p_2_8_11), .GIK(g_2_8_11), .GKJ(g_3_0_7), .GIJ(g_3_0_11));
GrayCell U31 (.PIK(p_1_4_5), .GIK(g_1_4_5), .GKJ(g_2_0_3), .GIJ(g_2_0_5));
GrayCell U32 (.PIK(p_1_8_9), .GIK(g_1_8_9), .GKJ(g_3_0_7), .GIJ(g_2_0_9));
GrayCell U33 (.PIK(p_1_12_13), .GIK(g_1_12_13), .GKJ(g_3_0_11), .GIJ(g_2_0_13));
GrayCell U34 (.PIK(p_0_2_2), .GIK(g_0_2_2), .GKJ(g_1_0_1), .GIJ(g_1_0_2));
GrayCell U35 (.PIK(p_0_4_4), .GIK(g_0_4_4), .GKJ(g_2_0_3), .GIJ(g_1_0_4));
GrayCell U36 (.PIK(p_0_6_6), .GIK(g_0_6_6), .GKJ(g_2_0_5), .GIJ(g_1_0_6));
GrayCell U37 (.PIK(p_0_8_8), .GIK(g_0_8_8), .GKJ(g_3_0_7), .GIJ(g_1_0_8));
GrayCell U38 (.PIK(p_0_10_10), .GIK(g_0_10_10), .GKJ(g_2_0_9), .GIJ(g_1_0_10));
GrayCell U39 (.PIK(p_0_12_12), .GIK(g_0_12_12), .GKJ(g_3_0_11), .GIJ(g_1_0_12));
GrayCell U40 (.PIK(p_0_14_14), .GIK(g_0_14_14), .GKJ(g_2_0_13), .GIJ(g_1_0_14));
assign S[16] = c[16];
assign c[0] = 1'b0;
assign c[10] = g_2_0_9;
assign c[11] = g_1_0_10;
assign c[12] = g_3_0_11;
assign c[13] = g_1_0_12;
assign c[14] = g_2_0_13;
assign c[15] = g_1_0_14;
assign c[16] = g_4_0_15;
assign c[1] = g_0_0_0;
assign c[2] = g_1_0_1;
assign c[3] = g_1_0_2;
assign c[4] = g_2_0_3;
assign c[5] = g_1_0_4;
assign c[6] = g_2_0_5;
assign c[7] = g_1_0_6;
assign c[8] = g_3_0_7;
assign c[9] = g_1_0_8;
xor UXOR0 (S[0], p_0_0_0, c[0]);
xor UXOR1 (S[1], p_0_1_1, c[1]);
xor UXOR10 (S[10], p_0_10_10, c[10]);
xor UXOR11 (S[11], p_0_11_11, c[11]);
xor UXOR12 (S[12], p_0_12_12, c[12]);
xor UXOR13 (S[13], p_0_13_13, c[13]);
xor UXOR14 (S[14], p_0_14_14, c[14]);
xor UXOR15 (S[15], p_0_15_15, c[15]);
xor UXOR2 (S[2], p_0_2_2, c[2]);
xor UXOR3 (S[3], p_0_3_3, c[3]);
xor UXOR4 (S[4], p_0_4_4, c[4]);
xor UXOR5 (S[5], p_0_5_5, c[5]);
xor UXOR6 (S[6], p_0_6_6, c[6]);
xor UXOR7 (S[7], p_0_7_7, c[7]);
xor UXOR8 (S[8], p_0_8_8, c[8]);
xor UXOR9 (S[9], p_0_9_9, c[9]);
endmodule