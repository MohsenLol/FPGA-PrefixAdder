library verilog;
use verilog.vl_types.all;
entity BrentKung64b_etb is
end BrentKung64b_etb;
