library verilog;
use verilog.vl_types.all;
entity KoggeStone16b_tb is
end KoggeStone16b_tb;
