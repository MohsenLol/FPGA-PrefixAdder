library verilog;
use verilog.vl_types.all;
entity BrentKung32b_tb is
end BrentKung32b_tb;
