library verilog;
use verilog.vl_types.all;
entity rippleCarry8b_tb is
end rippleCarry8b_tb;
