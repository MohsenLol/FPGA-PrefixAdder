library verilog;
use verilog.vl_types.all;
entity BrentKung16b_etb is
end BrentKung16b_etb;
