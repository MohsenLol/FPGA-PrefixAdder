library verilog;
use verilog.vl_types.all;
entity BrentKung16b_tb is
end BrentKung16b_tb;
