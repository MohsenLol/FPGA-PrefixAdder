library verilog;
use verilog.vl_types.all;
entity BrentKung8b_etb is
end BrentKung8b_etb;
