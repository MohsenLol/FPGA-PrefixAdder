module BrentKung8b (A, B, S);
input [7 : 0] A;
input [7 : 0] B;
output [8 : 0] S;
wire g_1_0_2, g_2_0_5, g_0_5_5, p_1_4_5, p_0_3_3, p_1_6_7, p_0_6_6, c [8 : 0], p_0_0_0, p_0_2_2, g_2_0_3, p_0_5_5, g_0_7_7, g_3_0_7, g_1_4_5, p_0_7_7, g_0_6_6, g_2_4_7, g_0_0_0, g_0_3_3, p_0_4_4, g_1_0_6, g_1_0_1, g_0_4_4, g_1_6_7, p_1_2_3, g_1_0_4, g_1_2_3, p_2_4_7, g_0_1_1, g_0_2_2, p_0_1_1;
BlackCell U10 (.PIK(p_0_7_7), .GIK(g_0_7_7), .GKJ(g_0_6_6), .PKJ(p_0_6_6),  .GIJ(g_1_6_7), .PIJ(p_1_6_7));
BlackCell U12 (.PIK(p_1_6_7), .GIK(g_1_6_7), .GKJ(g_1_4_5), .PKJ(p_1_4_5),  .GIJ(g_2_4_7), .PIJ(p_2_4_7));
BlackCell U8 (.PIK(p_0_3_3), .GIK(g_0_3_3), .GKJ(g_0_2_2), .PKJ(p_0_2_2),  .GIJ(g_1_2_3), .PIJ(p_1_2_3));
BlackCell U9 (.PIK(p_0_5_5), .GIK(g_0_5_5), .GKJ(g_0_4_4), .PKJ(p_0_4_4),  .GIJ(g_1_4_5), .PIJ(p_1_4_5));
GPCell UGP0 (.A(A[0]), .B(B[0]), .G(g_0_0_0), .P(p_0_0_0));
GPCell UGP1 (.A(A[1]), .B(B[1]), .G(g_0_1_1), .P(p_0_1_1));
GPCell UGP2 (.A(A[2]), .B(B[2]), .G(g_0_2_2), .P(p_0_2_2));
GPCell UGP3 (.A(A[3]), .B(B[3]), .G(g_0_3_3), .P(p_0_3_3));
GPCell UGP4 (.A(A[4]), .B(B[4]), .G(g_0_4_4), .P(p_0_4_4));
GPCell UGP5 (.A(A[5]), .B(B[5]), .G(g_0_5_5), .P(p_0_5_5));
GPCell UGP6 (.A(A[6]), .B(B[6]), .G(g_0_6_6), .P(p_0_6_6));
GPCell UGP7 (.A(A[7]), .B(B[7]), .G(g_0_7_7), .P(p_0_7_7));
GrayCell U11 (.PIK(p_1_2_3), .GIK(g_1_2_3), .GKJ(g_1_0_1), .GIJ(g_2_0_3));
GrayCell U13 (.PIK(p_2_4_7), .GIK(g_2_4_7), .GKJ(g_2_0_3), .GIJ(g_3_0_7));
GrayCell U14 (.PIK(p_1_4_5), .GIK(g_1_4_5), .GKJ(g_2_0_3), .GIJ(g_2_0_5));
GrayCell U15 (.PIK(p_0_2_2), .GIK(g_0_2_2), .GKJ(g_1_0_1), .GIJ(g_1_0_2));
GrayCell U16 (.PIK(p_0_4_4), .GIK(g_0_4_4), .GKJ(g_2_0_3), .GIJ(g_1_0_4));
GrayCell U17 (.PIK(p_0_6_6), .GIK(g_0_6_6), .GKJ(g_2_0_5), .GIJ(g_1_0_6));
GrayCell U7 (.PIK(p_0_1_1), .GIK(g_0_1_1), .GKJ(g_0_0_0), .GIJ(g_1_0_1));
assign S[8] = c[8];
assign c[0] = 1'b0;
assign c[1] = g_0_0_0;
assign c[2] = g_1_0_1;
assign c[3] = g_1_0_2;
assign c[4] = g_2_0_3;
assign c[5] = g_1_0_4;
assign c[6] = g_2_0_5;
assign c[7] = g_1_0_6;
assign c[8] = g_3_0_7;
xor UXOR0 (S[0], p_0_0_0, c[0]);
xor UXOR1 (S[1], p_0_1_1, c[1]);
xor UXOR2 (S[2], p_0_2_2, c[2]);
xor UXOR3 (S[3], p_0_3_3, c[3]);
xor UXOR4 (S[4], p_0_4_4, c[4]);
xor UXOR5 (S[5], p_0_5_5, c[5]);
xor UXOR6 (S[6], p_0_6_6, c[6]);
xor UXOR7 (S[7], p_0_7_7, c[7]);
endmodule