library verilog;
use verilog.vl_types.all;
entity LadnerFischer16b_tb is
end LadnerFischer16b_tb;
