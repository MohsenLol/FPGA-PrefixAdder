library verilog;
use verilog.vl_types.all;
entity BrentKung32b_rtb is
end BrentKung32b_rtb;
